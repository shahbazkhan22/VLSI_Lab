** Profile: "SCHEMATIC1-ResistiveLoad"  [ C:\Users\shahb\Documents\ResisitiveLoad-PSpiceFiles\SCHEMATIC1\ResistiveLoad.sim ] 

** Creating circuit file "ResistiveLoad.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../resisitiveload-pspicefiles/resisitiveload.lib" 
* From [PSPICE NETLIST] section of C:\Users\shahb\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 1.8 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
