** Profile: "SCHEMATIC1-PMos"  [ C:\Users\shahb\Documents\PMos-PSpiceFiles\SCHEMATIC1\PMos.sim ] 

** Creating circuit file "PMos.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../pmos-pspicefiles/pmos.lib" 
* From [PSPICE NETLIST] section of C:\Users\shahb\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V1 0 1.8 .01 
+ LIN V_V2 0 1.2 0.6 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
